library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity FSMClockUnit is
end FSMClockUnit;

architecture Behavioral of FSMClockUnit is

begin


end Behavioral;

