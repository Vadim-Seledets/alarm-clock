library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity AudioDriver is
	port (
		PlayEnable: in std_logic;
		CLK: in std_logic
	);
end AudioDriver;

architecture Behavioral of AudioDriver is

begin


end Behavioral;

